*
* NGSPICE simulation script
*

* forces current values to be saved
.options savecurrents

* include data for simulation when t<0
.INCLUDE data_sim.txt

.model P2model NPN(Bf=200, CJE=12pF, CJC=2pF)

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

print V(6)-V(8) > datav6v8.txt 
print V(6)-V(8) > dataic.txt
echo  "op_TAB"
print all
echo  "op_END"

quit
.endc

.end