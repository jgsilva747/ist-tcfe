*-------------------------------------------------------
* NGSPICE simulation script
* natural repsonse of circuit with boundary conditions v(6) and v(8) as computed in sim_t2_2.net

* forces current values to be saved
.options savecurrents

*resistors
.INCLUDE data_sim3.txt
.INCLUDE dataic.txt
*.ic v(6) = 8.573530 v(8) = 0 
*alterar para automatizar depois

.end 

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-6 20e-3

hardcopy trans.ps v(6) 
echo trans_FIG

quit
.endc
.end