T1 transient analysis

* NGSPICE simulation script
* BJT amp with feedback
*

* forces current values to be saved
.options savecurrents


*Resistors
R1 N1 N2 1.01658203395k
R2 N2 N3 2.08071598482k
R3 N2 N5 3.12527703197k
R4 0 N5 4.13615246449k
R5 N5 N6 3.04804224053k
R6 0 N4 2.06609096892k
R7 N7 N8 1.01589064139k

*Condensator
C N6 N8 1.02439571082u

*Independent Voltage and Current Sources
Vs N1 0 DC 0

Id N1 N2 DC 1.02439571082m

V3 N4 N7 DC 0

*Dependent Voltage and Current Sources

Gb N6 N3 N2 N5 7.30340439475m

Hc N5 N8 V3 8.13276803722k


.ic v(n6) = 9.707995e+00
.ic v(n8) = -6.12046e-01

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "****************"
echo  "Operating point"
echo "****************"
*print v-sweep
*print @R6[i]

*Tabela Principal

echo  "op2_TAB"
print all
echo  "op2_END"

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-3 20e-3

hardcopy naturaltrans.ps v(n6)
echo naturaltrans_FIG

.endc
.end